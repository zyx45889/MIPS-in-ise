`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:35:11 06/21/2020 
// Design Name: 
// Module Name:    SLL 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module SLL(
input [31:0]A,
input [5:0]B,
output [31:0]C
    );
//uncompleted
assign C=A;

endmodule