`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:32:17 04/23/2020 
// Design Name: 
// Module Name:    SRL 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module SRL(
input [31:0]A,
input [5:0]B,
output [31:0]C
    );
//uncompleted
assign C=A;

endmodule
